'00000000000000000000000000000000'001000 0 101',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 101 101',
'00000000000000000000000000000000'00000000000000000000000000000000'001000 0 101',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 110 101',
'00000000000000000000000000000000'00000000000000000000000000000000'101011 0 101',
'00000000000000000000000000000000'00000000000000000000000000000000'100011 0 111',
'00000000000000000000000000000000'00000000000000000000000000000000'001000 0 100',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 100 101',
'00000000000000000000000000000000'00000000000000000000000000000000'001100 100 100',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 111 11',
'00000000000000000000000000000000'00000000000000000000000000000000'001101 101 101',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 101 111',
'00000000000000000000000000000000'00000000000000000000000000000000'001000 0 1',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 111 1',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 111 1',
'00000000000000000000000000000000'00000000000000000000000000000000'001010 111 11',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 1 1',
'00000000000000000000000000000000'00000000000000000000000000000000'000000 111 111',
'00000000000000000000000000000000'00000000000000000000000000000000'000100 0 11',
'00000000000000000000000000000000'00000000000000000000000000000000'00000000000000000000000000000000'00000000000000000000000000000000'00000000000000000000000000000000'001000 0 10',
'00000000000000000000000000000000'00000000000000000000000000000000'000101 111 10',
'001000 111 111',
'001000 111 111',
'00000000000000000000000000000000(others => '1'),
others => (others => '0')